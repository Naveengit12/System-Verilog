// INTERFACE

interface and_gate;
  logic a,b;
  logic y;
endinterface
