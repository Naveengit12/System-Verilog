
module four_state_datatype;
  wire a;
  reg b;
  logic c;
  time d;
  integer e;
  real f;

  initial begin
    $display("a=%b, b=%b, c=%b, d=%0d, e=%d,f=%0d", a, b, c, d, e, f);
  end
endmodule
