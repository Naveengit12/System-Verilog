module four_state_datatype;
  wire a;
  reg b;
  logic c;
  time d;
  integer e;
  initial begin
    $display("a=%d, b=%d, c=%d, d=%0d, e=%d", a, b, c, d, e);
  end
endmodule
