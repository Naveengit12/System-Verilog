module four_state_datatype;
  wire a;
  reg b;
  logic c;
  time d;
  integer e;
  real f;
  
  initial begin
    $display("a=%d, b=%d, c=%d, d=%0d, e=%d, f=%d", a, b, c, d, e, f);
  end
endmodule
