module two_state_datatype;
int a;
shortint b;
longint c;
real f;
bit e;
byte d;

initial begin
$display(" a=%b, b=%b, c=%b, d=%b, e=%b, f=%f", a,b,c,d,e,f);
end
endmodule
