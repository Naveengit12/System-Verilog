// DESIGN PART

module andgate(and_gate Ag);
  assign Ag.y = Ag.a & Ag.b;
endmodule
