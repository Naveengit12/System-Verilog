module two_state_datatype;
int a;
shortint b;
longint c;
bit e;
byte d;

initial begin
$display(" a=%b, b=%b, c=%b, d=%b, e=%b", a,b,c,d,e,f);
end
endmodule
