// INTERFACE

interface full_adder;
  logic a,b,C_in;
  logic sum,C_out;
endinterface
