/*write a code for queue array with 4 elements... insert 1in the 1st index.. delete element in
3rd index... insert 9 as the last element... shuffle, reverse the elements  */
