/*write a code for dynamic array... give the value of array using foreach.. display the size..shuffle the array elements.../*

