// -------------------FORK JOIN---------------------------
module fork_join;
  
  initial begin
    fork
      begin
        $display("A is going GYM at time = %0t",$time);
        #15;
        $display("A is reached GYM at time = %0t",$time);
      end
      
      begin
        $display("B is doing workout at time = %0t",$time);
        #20;
        $display("B is completed workout at time = %0t",$time);
      end
      
      begin
        $display("A is started workout at time = %0t",$time);
        #20;
        $display("A is completed workout at time = %0t",$time);
      end
    join
  end
endmodule




// output
// # run -all
// # A is going GYM at time = 0
// # B is doing workout at time = 0
// # A is started workout at time = 0
// # A is reached GYM at time = 15
// # B is completed workout at time = 20
// # A is completed workout at time = 20
// # exit
