/*Create a typdef Instr_t of struct for the instruction and then declare the memory as array of
Instr_t */

